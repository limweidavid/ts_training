`define INPUT_SKEW 1
`define OUTPUT_SKEW 1