///////////////////////////////////////////////////////////////////////////
//
// File name         : 
// Author            : Shamaim
// Creation Date     : January 1st, 2024
//
// No portions of this material may be reproduced in any form without
// the written permission of Thundersoft
//
// No portions of this material may be reproduced in any form without
// the written permission of Thundersoft
//
// Description : 
//
///////////////////////////////////////////////////////////////////////////

`include "uvm_macros.svh"
package fifo_uvc_package;
  import uvm_pkg::*;

  `include "env/uvc/fifo/sequence_item.sv"
  `include "env/uvc/fifo/sequencer.sv"
  `include "env/uvc/fifo/driver.sv"
  `include "env/uvc/fifo/monitor.sv"
  `include "env/uvc/fifo/agent.sv"
endpackage